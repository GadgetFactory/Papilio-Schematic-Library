----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:01:17 11/27/2013 
-- Design Name: 
-- Module Name:    MISC_zpuino_sa_splitter4 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MISC_zpuino_sa_splitter4 is
    Port ( in1 : in  STD_LOGIC;
           out1 : out  STD_LOGIC;
			  out2 : out  STD_LOGIC;
			  out3 : out  STD_LOGIC;
           out4 : out  STD_LOGIC);
end MISC_zpuino_sa_splitter4;

architecture Behavioral of MISC_zpuino_sa_splitter4 is

begin
out1 <= in1;
out2 <= in1;
out3 <= in1;
out4 <= in1;

end Behavioral;

